


module fibonacci_top
